`define NONE 0

// Operations
`define PUSH    1
`define POP     2
`define REPLACE 3

// Status
`define UNDERFLOW 1
`define EMPTY     2
`define FULL      3

// Errors
`define OVERFLOW 2
